module TB;
    
endmodule
